-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Wednesday, May 21, 2014 07:07:16 SE Asia Standard Time

